//
// coding convention Dudy October 2020
// (c) Technion IIT, Department of Electrical Engineering 2019 
// generating a number bitmap 



module diamondsMatrices	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] pixelX,// offset from top left  position 
					input 	logic	[10:0] pixelY,
					input		logic	collision, //input that the pixel is within a bracket 
					input 	logic	[3:0] level, // digit to display
					
					
					output	logic	drawingRequest //output that the pixel should be dispalyed 
					//output	logic	[7:0]		RGBout
);
// generating a smily bitmap 

//parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 

//logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {

//RGBout <= object_colors[(pixelY - topLeftY)][(pixelX - topLeftX)];

//middle is length of each matrix ///rhs is size of row

logic [0:7-1] [0:15-1] [0:20-1] objects_position;
logic [0:7-1] [0:15-1] [0:20-1] objects_position0 = {

//level1
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000010000000000,
20'b	00000000000000000000,
20'b	00000111010101000000,
20'b	00000000000000010000,
20'b	00110000000100000000,
20'b	00000000010010100000,
20'b	00000000100000000000,
20'b	00000001000000000000,
20'b	00000000000000100000,
20'b	00011000000000000000,
20'b	00000011000000000000,
20'b	00000000000000000000,




},

//level2
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000110000000000000,
20'b	00000000000000000000,
20'b	00000000001010000000,
20'b	00000000000000000000,
20'b	00000000001110000000,
20'b	00000000000100000000,
20'b	00001000000000000000,
20'b	00000001000000000000,
20'b	00001100000000000000,
20'b	00000000000000000000,
20'b	00011001100000000000,
20'b	00000000000000000000,
},

//level3
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000011100001000000,
20'b	00001100000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00001111000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00100000000000111000,
20'b	00000000010000001100,
20'b	00000000000000000000,


},

//level4
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000011100,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000100000000000,
20'b	01111000000000000000,
20'b	00000000000000000000,
20'b	00010011111000000000,
20'b	00000000000000000000,
},


//level5
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00011111000011111000,
20'b	00011111100111110000,
20'b	00001111111111100000,
20'b	00000111111111100000,
20'b	00000011111110000000,
20'b	00000011000111000000,
20'b	00000001111111100000,
20'b	00001111111111110000,
20'b	00011111100111111000,
20'b	00011110000011111000,
20'b	00011100000000111000,
20'b	00000000000000000000,
},

//level6
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000010000000000000,
20'b	00001000101001111000,
20'b	00000000001001111000,
20'b	00010000000001111000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00010000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000111000,
20'b	00111000001111000000,
20'b	00000000000000000000,
},

//level7 -MAZE
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	01110000010111000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	01100000000000000000,
20'b	00001100000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000011100000000000,
20'b	00000000000000000000,
20'b	00000000000000111100,
20'b	00001110000000100100,
20'b	00000000000000000000,
},

};


// pipeline (ff) to get the pixel color from the array 	 

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
		objects_position <=objects_position0;
	end
	else begin
			//drawingRequest <= (objects_position[digit][offsetY][offsetX]) && (InsideRectangle == 1'b1 );	//get value from bitmap  
		if (objects_position[level][pixelY >> 5][pixelX >> 5]) begin /*&& (InsideRectangle == 1'b1*/ 
			drawingRequest <= 1;
		if (collision)
			objects_position[level][pixelY >> 5][pixelX >> 5] <=0;
		end
		else
			drawingRequest <= 0;
	end 
end

//assign RGBout = digit_color ; // this is a fixed color 

endmodule