//
// coding convention Dudy October 2020
// (c) Technion IIT, Department of Electrical Engineering 2019 
// generating a number bitmap 



module minesMatrices	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] pixelX,// offset from top left  position 
					input 	logic	[10:0] pixelY,
					input		logic	collision, //input that the pixel is within a bracket 
					input 	logic	[3:0] level, // digit to display
					
					
					output	logic	drawingRequest //output that the pixel should be dispalyed 
					//output	logic	[7:0]		RGBout
);
// generating a smily bitmap 

//parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 

//logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {

//RGBout <= object_colors[(pixelY - topLeftY)][(pixelX - topLeftX)];

//middle is length of each matrix ///rhs is size of row
logic [0:7-1] [0:15-1] [0:20-1] objects_position;

//7 levels , 15 rows to represent y, 20 columns to represent x
logic [0:7-1] [0:15-1] [0:20-1] objects_position0= {

//level1
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000001000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000010000,
20'b	00000000010000000000,
20'b	00000000000000000000,




},

//level2
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000100000000,
20'b	00000000000000000000,
20'b	00000000000100000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000010000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000110000000000000,
20'b	00000000000000000000,
},

//level3
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000100000,
20'b	00000000000000000000,
20'b	01100000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00010000000000000000,
20'b	00000000000001000000,
20'b	00000000000000000000,


},

//level4
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000100000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000001100000000,
20'b	00100000000000000000,
20'b	00000000000000000000,
},


//level5
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00110000000000000000,
20'b	00000000000000000000,
20'b	00000000000000001100,
20'b	00000000111000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000001100000000000,
20'b	00000000000000000000,
},

//level6
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000100,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	01000000110000011000,
20'b	00000000000000000000,
},

//level7 -MAZE
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000010000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	01000000000000000000,
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	00000001000000000000,
20'b	00000000000000011000,
20'b	00000000000000000000,
},

};


// pipeline (ff) to get the pixel color from the array 	 

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
		objects_position <=objects_position0;
		end
	else begin
			//drawingRequest <= (objects_position[digit][offsetY][offsetX]) && (InsideRectangle == 1'b1 );	//get value from bitmap  
		if (objects_position[level][pixelY >> 5][pixelX >> 5]) begin /*&& (InsideRectangle == 1'b1*/ 
			drawingRequest <= 1;
		if (collision)
			objects_position[level][pixelY >> 5][pixelX >> 5] <=0;
		end
		else
			drawingRequest <= 0;
	end 
end

//assign RGBout = digit_color ; // this is a fixed color 

endmodule