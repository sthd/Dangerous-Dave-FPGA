//
// coding convention Dudy October 2020
// (c) Technion IIT, Department of Electrical Engineering 2019 
// generating a number bitmap 



module blocksMatrices	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] pixelX,// offset from top left  position 
					input 	logic	[10:0] pixelY,
					input		logic	collision, //input that the pixel is within a bracket 
					input 	logic	[3:0] level, // digit to display
					
					
					output	logic	drawingRequest //output that the pixel should be dispalyed 
					//output	logic	[7:0]		RGBout
);
// generating a smily bitmap 

//parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 

//logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {

//RGBout <= object_colors[(pixelY - topLeftY)][(pixelX - topLeftX)];

//middle is length of each matrix ///rhs is size of row
logic [0:7-1] [0:15-1] [0:20-1] objects_position;

logic [0:7-1] [0:15-1] [0:20-1] objects_position0 = {

//level1
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000111000000000001,
20'b	10000000000000110001,
20'b	10110000011110000001,
20'b	10000001000000000001,
20'b	10000100000000000001,
20'b	10011000000000000001,
20'b	10000000000011110001,
20'b	10000001100000000001,
20'b	10000010000110100001,
20'b	10001000000001001001,
20'b	11111111111111111111,
},

//level2
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10110000001110001001,
20'b	10000110000000010001,
20'b	10000000111111000001,
20'b	10011110000000000001,
20'b	10000000001010010101,
20'b	10000000011111000001,
20'b	10011110000000000001,
20'b	10000000000111111101,
20'b	10011111110000000001,
20'b	10000000000000000001,
20'b	11111111111111111111,
},

//level3
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000000000111110001,
20'b	10011110000000000001,
20'b	10000000000001100001,
20'b	10000000011100000001,
20'b	10011000000000011001,
20'b	10000010100000111111,
20'b	10011111111000000001,
20'b	10100000000011100001,
20'b	10001110111000000001,
20'b	10111000000000000001,
20'b	11111111111111111111,

},

//level4
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000001111111000001,
20'b	10000011111111110001,
20'b	10001111111111110001,
20'b	10011111111111000001,
20'b	10011111100111001001,
20'b	10011110000011001001,
20'b	10011100000011001001,
20'b	10000000000001001101,
20'b	10000000110001001001,
20'b	10000011110001001001,
20'b	10000000000001001001,
20'b	11111111111111111111,
},


//level5
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000110000000011111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000001111000000001,
20'b	10000000000000000001,
20'b	11111111111111111111,
},

//level6
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10011110100110000001,
20'b	10000000101000000001,
20'b	10111000101001100001,
20'b	10000011101000001101,
20'b	10000000101000011001,
20'b	10011000101001100001,
20'b	10000000000000000001,
20'b	11110011111110000101,
20'b	10000000000000000001,
20'b	11111111111111111111,
},

//level7 -MAZE
{
20'b	00000000000000000000,
20'b	00000000000000000000,
20'b	11111111111111111111,
20'b	10000000001000000101,
20'b	10110111010100101001,
20'b	10110010001010001011,
20'b	10001100000111000001,
20'b	10000001011000110111,
20'b	10011100010011000001,
20'b	10000001111000001111,
20'b	10011100000011100001,
20'b	10000001100110000001,
20'b	10011010001000000001,
20'b	10000000010000000001,
20'b	11111111111111111111,
},

};

/*
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;

//4 levels , 15 rows to represent y, 20 columns to represent x
objects_position <
	end
end
*/

// pipeline (ff) to get the pixel color from the array 	 

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
		objects_position <=objects_position0;
	end
	else begin
			//drawingRequest <= (objects_position[digit][offsetY][offsetX]) && (InsideRectangle == 1'b1 );	//get value from bitmap  
		if (objects_position[level][pixelY >> 5][pixelX >> 5]) begin /*&& (InsideRectangle == 1'b1*/ 
			drawingRequest <= 1;
		if (collision)
			objects_position[level][pixelY >> 5][pixelX >> 5] <=0;
		end
		else
			drawingRequest <= 0;
	end 
end

//assign RGBout = digit_color ; // this is a fixed color 

endmodule